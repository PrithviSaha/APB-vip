//`include "defines.svh"
class apb_driver extends uvm_driver #(apb_sequence_item);
  `uvm_component_utils(apb_driver)

  virtual apb_if vif;
  
 // uvm_analysis_port #(apb_sequence_item) item_collected_port;   //port for coverage
    
  function new (string name = "apb_driver", uvm_component parent );
    super.new(name, parent);
   // item_collected_port = new("item_collected_port", this);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    if(!uvm_config_db#(virtual apb_if)::get(this, "", "vif", vif))
       `uvm_fatal("NO_VIF",{"virtual interface must be set for: ",get_full_name(),".vif"});

  endfunction
  
  task send_to_interface();
    vif.drv_cb.PRESETn <= req.PRESETn;
    vif.drv_cb.transfer <= req.transfer;
    vif.drv_cb.READ_WRITE <= req.READ_WRITE;
    vif.drv_cb.apb_read_paddr <= req.apb_read_paddr;
    vif.drv_cb.apb_write_paddr <= req.apb_write_paddr;
    vif.drv_cb.apb_write_data <= req.apb_write_data;
  endtask

  task drive();
    send_to_interface();
    repeat(2) @(posedge vif.PCLK)
  endtask

  task run_phase(uvm_phase phase);
    repeat(3) @(posedge vif.PCLK);
    forever begin
      seq_item_port.get_next_item(req);
      drive();
      seq_item_port.item_done();
    end
  endtask   

endclass
