`define DATA_WIDTH 8;
`define ADDR_WISTH 9;

