package alp_pkg;
  `include "apb_sequence_item.sv"
  `include "apb_sequence.sv"
  `include "apb_sequencer.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_active_agent.sv"
  `include "apb_passive_agent.sv"
  `include "apb_input_monitor.sv"
   `include "apb_input_monitor.sv"
  `include "apb_scoreboard.sv"
 `include "apb_coverage.sv"
  `include "apb_environment.sv"
  `include "apb_test.sv"
  `include "defines.svh"
endpackage
