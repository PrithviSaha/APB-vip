`define ADDR_WIDTH 9
`define WIDTH 8
